library ieee;
use ieee.std_logic_1164.all;
use ieee.numeric_std.all;

package Synthesis_definitions_pack is
	constant maximum_multiplier_width : integer := 16; -- 18 maximo para la spartan6, para la kintex7 es 25x18
end package;

package body Synthesis_definitions_pack is
end package body;